module firpga (              
	input                     sys_clk,
	input                     sys_rst,
	//////////////
	//audio part//
	//////////////
	//WM978 interface
	input                     aud_bclk,   //bit clk
	input                     aud_lrc,    //synchronize signal
	input                     aud_adcdat, //audio_input
	input                     key0,
	output                    aud_mclk,   //main clk signal for WM8978,generated by pll ip core
	output                    aud_dacdat,  //audio output
	//control interface
	output                    aud_scl,    //WM8978 audio IIC clock signal
	inout                     aud_sda,    //WM8978 audio IIC data signal
	
	////////////
	//fft part//
	////////////
	
	////////////
	//lcd part//
	////////////
	output                    lcd_hs,
	output                    lcd_vs,
	output                    lcd_de,
	output      [15:0]        lcd_rgb,
	output                    lcd_bl,
	output                    lcd_rst,
	output                    lcd_pclk
);

//parameter define


//reg define

//wire define
wire    [15:0]      adc_data;   //audio data sampled by FPGA
wire    [15:0]      overdrive_data;   //audio output form the fir filter
wire                rx_done;    //an output from the audio interface
//signals connecting the fft module and the lcd_top module
wire                fft_valid;  //output of the fft module data_valid
//wire                fir_valid;  //output of the fir module data_valid
wire                fft_sop;
wire                fft_eop;
wire    [15:0]      fft_data;   //output of the fft module data_modulus
wire    [15:0]      audio_data_out; //the data going to the wm8978 input port

//************************************************************************************
//                 main code
//************************************************************************************
assign audio_data_out = key0?overdrive_data:adc_data; //if press the button key0 then output is filtered data
//the audio part
//the pll module is just to generate a 12MHz signal and to be the main clock signal of the chip
pll_clk u_pll_clk(
    .areset             (~sys_rst  ),   
    .inclk0             (sys_clk   ),   
    .c0                 (aud_mclk  )    //the output to be the clock of the chip
);

//WM8978 control
wm8978_ctrl u_wm8978_ctrl(
    .clk                (sys_clk    ),  
    .rst_n              (sys_rst    ),  

    .aud_bclk           (aud_bclk   ),  //clk signal coming from the chip, control the data transmission
    .aud_lrc            (aud_lrc    ),  //synchronization signal
    .aud_adcdat         (aud_adcdat ),  //data transmission
    .aud_dacdat         (aud_dacdat ),  
    
    .aud_scl            (aud_scl    ),  //scl signal of IIC
    .aud_sda            (aud_sda    ),  //SDA signal of IIC
    
    .adc_data           (adc_data   ),  
    .dac_data           (audio_data_out   ),  /////////need to be changed to fir_data//////////////////////////
    .rx_done            (rx_done),             
    .tx_done            ()              
);


//the fft_part
fft_top u_fft_top(
	.sys_clk             (sys_clk),
	.sys_rst             (sys_rst),
	
	.audio_clk           (aud_bclk),
	.audio_data          (audio_data_out),
	.audio_valid         (rx_done),
	
	.data_sop            (fft_sop),
	.data_eop            (fft_eop),
	.data_valid          (fft_valid),
	.data_modulus        (fft_data)
);


//the LCD part
lcd_top u_lcd_top(
	.sys_clk             (sys_clk),
	.sys_rst             (sys_rst),
	//signal coming from the fft module
	.fft_data            (fft_data),
	.fft_sop             (fft_sop),
	.fft_eop             (fft_eop),
	.fft_valid           (fft_valid),
	//signal going to the lcd display
	.lcd_bl              (lcd_bl),
	.lcd_de              (lcd_de),
	.lcd_rgb             (lcd_rgb),
	.lcd_vs              (lcd_vs),
	.lcd_hs              (lcd_hs),
	.lcd_rst             (lcd_rst),
	.lcd_pclk            (lcd_pclk)
);

//fir filter module, get data from the receiver and do filtering
overdrive u_overdrive(
	 .clk            (aud_bclk),
	 .reset          (sys_rst),
	 //audio input 
	 .clk_enable     (rx_done),
	 .overdrive_in       (adc_data),
	 //output signals
	 .overdrive_out      (overdrive_data),

);
endmodule
