/*
30/6/2021
created by ALIENTEK. Co
modified by Zyy Zhou (22670661)
this file is to realize an audio encoder chip and let the data
go through the FPGA inside. then let the audio data go back to 
the wm8978 chip without processing the signal
*/
module audio_speak (
	input                     sys_clk,
	input                     sys_rst,
	//WM978 interface
	input                     aud_bclk,   //bit clk
	input                     aud_lrc,    //synchronize signal
	input                     aud_adcdat, //audio_input
	output                    aud_mclk,   //main clk signal for WM8978,generated by pll ip core
	output                    aud_dacdat,  //audio output
	//control interface
	output                    aud_scl,    //WM8978 audio IIC clock signal
	inout                     aud_sda    //WM8978 audio IIC data signal
);

//parameter define

//reg define

//wire define
wire    [31:0]      adc_data;   //audio data sampled by FPGA

//***********************************************************************
//                       main code
//***********************************************************************

//the pll module is just to generate a 12MHz signal and to be the main clock signal of the chip
pll_clk u_pll_clk(
    .areset             (~sys_rst  ),   
    .inclk0             (sys_clk   ),   
    .c0                 (aud_mclk  )    //the output to be the clock of the chip
);

//WM8978 control
wm8978_ctrl u_wm8978_ctrl(
    .clk                (sys_clk    ),  
    .rst_n              (sys_rst    ),  

    .aud_bclk           (aud_bclk   ),  //clk signal coming from the chip, control the data transmission
    .aud_lrc            (aud_lrc    ),  //synchronization signal
    .aud_adcdat         (aud_adcdat ),  //data transmission
    .aud_dacdat         (aud_dacdat ),  
    
    .aud_scl            (aud_scl    ),  //scl signal of IIC
    .aud_sda            (aud_sda    ),  //SDA signal of IIC
    
    .adc_data           (adc_data   ),  
    .dac_data           (adc_data   ),  
    .rx_done            (),             
    .tx_done            ()              
);

endmodule 





