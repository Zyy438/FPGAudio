module fftpga (              
	input                     sys_clk,
	input                     sys_rst,
	//////////////
	//audio part//
	//////////////
	//WM978 interface
	input                     aud_bclk,   //bit clk
	input                     aud_lrc,    //synchronize signal
	input                     aud_adcdat, //audio_input
	output                    aud_mclk,   //main clk signal for WM8978,generated by pll ip core
	output                    aud_dacdat,  //audio output
	//control interface
	output                    aud_scl,    //WM8978 audio IIC clock signal
	inout                     aud_sda,    //WM8978 audio IIC data signal
	
	////////////
	//fft part//
	////////////
	
	////////////
	//lcd part//
	////////////
	output                    lcd_hs,
	output                    lcd_vs,
	output                    lcd_de,
	output      [15:0]        lcd_rgb,
	output                    lcd_bl,
	output                    lcd_rst,
	output                    lcd_pclk
);

//parameter define


//reg define

//wire define
wire    [31:0]      adc_data;   //audio data sampled by FPGA
wire                rx_done;    //an output from the audio interface
//signals connecting the fft module and the lcd_top module
wire                fft_valid;  //output of the fft module data_valid
wire                fft_sop;
wire                fft_eop;
wire    [15:0]      fft_data;   //output of the fft module data_modulus


//************************************************************************************
//                 main code
//************************************************************************************
//the audio part
//the pll module is just to generate a 12MHz signal and to be the main clock signal of the chip
pll_clk u_pll_clk(
    .areset             (~sys_rst  ),   
    .inclk0             (sys_clk   ),   
    .c0                 (aud_mclk  )    //the output to be the clock of the chip
);

//WM8978 control
wm8978_ctrl u_wm8978_ctrl(
    .clk                (sys_clk    ),  
    .rst_n              (sys_rst    ),  

    .aud_bclk           (aud_bclk   ),  //clk signal coming from the chip, control the data transmission
    .aud_lrc            (aud_lrc    ),  //synchronization signal
    .aud_adcdat         (aud_adcdat ),  //data transmission
    .aud_dacdat         (aud_dacdat ),  
    
    .aud_scl            (aud_scl    ),  //scl signal of IIC
    .aud_sda            (aud_sda    ),  //SDA signal of IIC
    
    .adc_data           (adc_data   ),  
    .dac_data           (adc_data   ),  
    .rx_done            (rx_done),             
    .tx_done            ()              
);


//the fft_part
fft_top u_fft_top(
	.sys_clk             (sys_clk),
	.sys_rst             (sys_rst),
	
	.audio_clk           (aud_bclk),
	.audio_data          (adc_data),
	.audio_valid         (rx_done),
	
	.data_sop            (fft_sop),
	.data_eop            (fft_eop),
	.data_valid          (fft_valid),
	.data_modulus        (fft_data)
);


//the LCD part
lcd_top u_lcd_top(
	.sys_clk             (sys_clk),
	.sys_rst             (sys_rst),
	//signal coming from the fft module
	.fft_data            (fft_data),
	.fft_sop             (fft_sop),
	.fft_eop             (fft_eop),
	.fft_valid           (fft_valid),
	//signal going to the lcd display
	.lcd_bl              (lcd_bl),
	.lcd_de              (lcd_de),
	.lcd_rgb             (lcd_rgb),
	.lcd_vs              (lcd_vs),
	.lcd_hs              (lcd_hs),
	.lcd_rst             (lcd_rst),
	.lcd_pclk            (lcd_pclk)
);


endmodule
